//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   File Name   : WD.v
//   Module Name : WD
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module WD(
    // Input signals
    clk,
    rst_n,
    in_valid,
    keyboard,
    answer,
    weight,
    match_target,
    // Output signals
    out_valid,
    result,
    out_value
);

// ===============================================================
// Input & Output Declaration
// ===============================================================
input clk, rst_n, in_valid;
input [4:0] keyboard, answer;
input [3:0] weight;
input [2:0] match_target;
output reg out_valid;
output reg [4:0]  result;
output reg [10:0] out_value;

// ===============================================================
// Parameters & Integer Declaration
// ===============================================================
parameter STATE_IDLE = 5'd0; // Initialization, store 1st input value when in_valid is triggered
parameter STATE_INPUT = 5'd1; // Store 2nd - 8th input value
parameter STATE_REORDER = 5'd2; // Reorder input along answer to iterate permutations
parameter STATE_5A0B = 5'd3; // 17 different types of NANB, 1 permutations
parameter STATE_4A0B = 5'd4; // 15 permutations
parameter STATE_3A2B = 5'd5; // 10 permutations
parameter STATE_3A1B = 5'd6; // 60 permutations
parameter STATE_3A0B = 5'd7; // 60 permutations
parameter STATE_2A3B = 5'd8; // 20 permutations
parameter STATE_2A2B = 5'd9; // 270 permutations
parameter STATE_2A1B = 5'd10; // 360 permutations
parameter STATE_2A0B = 5'd11; // 60 permutations
parameter STATE_1A4B = 5'd12; // 45 permutations
parameter STATE_1A3B = 5'd13; // 660 permutations
parameter STATE_1A2B = 5'd14; // 1260 permutations
parameter STATE_1A1B = 5'd15; // 360 permutations
parameter STATE_0A5B = 5'd16; // 44 permutations
parameter STATE_0A4B = 5'd17; // 795 permutations
parameter STATE_0A3B = 5'd18; // 1920 permutations
parameter STATE_0A2B = 5'd19; // 780 permutations
parameter STATE_OUTPUT = 5'd20;

// ===============================================================
// Wire & Reg Declaration
// ===============================================================
reg [4:0] current_state, next_state;
reg [10:0] cnt; // counter used for counting cycles to update FSM
reg [4:0] keyboard_arr[7:0]; // storing keyboard sequence
reg [4:0] reorder_arr[7:0]; // storing reorder sequence along answer sequence (may be combined with keyboard_arr TBD)
reg [4:0] answer_arr[4:0]; // storing answer sequence
reg [3:0] weight_arr[4:0]; // storing weight sequence
reg [2:0] match_target_arr[1:0]; // {A,B}
reg [4:0] perm_arr[4:0]; // iterating permutation candidates
reg [4:0] prev_perm_arr[4:0]; // temp saving for updating result in following cycles
reg [4:0] result_arr[4:0]; // storing result sequence
reg [13:0] weighted_sum, weighted_sum_2; // calculating weighted sum & corner case 1 weighted sum
reg [13:0] max_weighted_sum, max_weighted_sum_2; // storing max weighted sum
reg [24:0] bwnc; // calculating bitwise not concatenation for corner case 2
reg [24:0] max_bwnc; // storing max bwnc

genvar vi;
integer ii;

// ===============================================================
// DESIGN
// ===============================================================


// ===============================================================
// Finite State Machine
// ===============================================================
// Current State
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) current_state <= STATE_IDLE;
    else        current_state <= next_state;
end

// Next State
always @(*) begin
    if (!rst_n) next_state = STATE_IDLE;
    else begin
        case (current_state)
            STATE_IDLE: begin
                if (in_valid) next_state = STATE_INPUT;
                else next_state = current_state;
            end
            STATE_INPUT: begin // processing (cnt+2)th value
                if (cnt==6) next_state = STATE_REORDER;
                else next_state = current_state;
            end
            STATE_REORDER: begin 
                if (cnt==11'd25) begin // cnt+1 cycles required 
                    case ({match_target_arr[0],match_target_arr[1]})
                        {3'd5,3'd0}: next_state = STATE_5A0B;
                        {3'd4,3'd0}: next_state = STATE_4A0B;
                        {3'd3,3'd2}: next_state = STATE_3A2B;
                        {3'd3,3'd1}: next_state = STATE_3A1B;
                        {3'd3,3'd0}: next_state = STATE_3A0B;
                        {3'd2,3'd3}: next_state = STATE_2A3B;
                        {3'd2,3'd2}: next_state = STATE_2A2B;
                        {3'd2,3'd1}: next_state = STATE_2A1B;
                        {3'd2,3'd0}: next_state = STATE_2A0B;
                        {3'd1,3'd4}: next_state = STATE_1A4B;
                        {3'd1,3'd3}: next_state = STATE_1A3B;
                        {3'd1,3'd2}: next_state = STATE_1A2B;
                        {3'd1,3'd1}: next_state = STATE_1A1B;
                        {3'd0,3'd5}: next_state = STATE_0A5B;
                        {3'd0,3'd4}: next_state = STATE_0A4B;
                        {3'd0,3'd3}: next_state = STATE_0A3B;
                        {3'd0,3'd2}: next_state = STATE_0A2B;
                        default: next_state = current_state;
                    endcase
                end
                else next_state = current_state;
            end
            // Idea:
            // 0th cycle: read 1st permutation
            // 1st cycle: read 2nd permutation, calculate 1st weighted sum
            // 2nd cycle: read 3rd permutation, calculate 2nd weighted sum, update 1st result
            // 3rd cycle: read 4th permutation, calculate 3rd weighted sum, update 2nd result
            // ...... (requires no. of permutation + 2 cycles in total)
            STATE_5A0B: begin if (cnt==11'd2) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_4A0B: begin if (cnt==11'd16) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_3A2B: begin if (cnt==11'd11) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_3A1B: begin if (cnt==11'd61) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_3A0B: begin if (cnt==11'd61) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_2A2B: begin if (cnt==11'd271) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_2A3B: begin if (cnt==11'd21) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_2A1B: begin if (cnt==11'd361) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_2A0B: begin if (cnt==11'd61) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_1A4B: begin if (cnt==11'd46) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_1A3B: begin if (cnt==11'd661) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_1A2B: begin if (cnt==11'd1261) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_1A1B: begin if (cnt==11'd361) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_0A4B: begin if (cnt==11'd796) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_0A5B: begin if (cnt==11'd45) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_0A3B: begin if (cnt==11'd1921) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_0A2B: begin if (cnt==11'd781) next_state = STATE_OUTPUT; else next_state = current_state; end
            STATE_OUTPUT: begin if (cnt==11'd4) next_state = STATE_IDLE; else next_state = current_state; end // cnt+1 cycles required 
            default: next_state = current_state;
        endcase
    end
end

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) cnt <= 11'd0;
    else 
        case (current_state) // could use a larger case statement to share the adder resource TBD
            STATE_IDLE: cnt <= 11'd0;
            STATE_INPUT: if (cnt==11'd6) cnt <= 0; else cnt <= cnt + 1;
            STATE_REORDER: if (cnt==11'd25) cnt <= 0; else cnt <= cnt + 1;
            STATE_5A0B: if (cnt==11'd2) cnt <= 0; else cnt <= cnt + 1;
            STATE_4A0B: if (cnt==11'd16) cnt <= 0; else cnt <= cnt + 1;
            STATE_3A2B: if (cnt==11'd11) cnt <= 0; else cnt <= cnt + 1;
            STATE_3A1B: if (cnt==11'd61) cnt <= 0; else cnt <= cnt + 1;
            STATE_3A0B: if (cnt==11'd61) cnt <= 0; else cnt <= cnt + 1;
            STATE_2A2B: if (cnt==11'd271) cnt <= 0; else cnt <= cnt + 1;
            STATE_2A3B: if (cnt==11'd21) cnt <= 0; else cnt <= cnt + 1;
            STATE_2A1B: if (cnt==11'd361) cnt <= 0; else cnt <= cnt + 1;
            STATE_2A0B: if (cnt==11'd61) cnt <= 0; else cnt <= cnt + 1;
            STATE_1A4B: if (cnt==11'd46) cnt <= 0; else cnt <= cnt + 1;
            STATE_1A3B: if (cnt==11'd661) cnt <= 0; else cnt <= cnt + 1;
            STATE_1A2B: if (cnt==11'd1261) cnt <= 0; else cnt <= cnt + 1;
            STATE_1A1B: if (cnt==11'd361) cnt <= 0; else cnt <= cnt + 1;
            STATE_0A4B: if (cnt==11'd796) cnt <= 0; else cnt <= cnt + 1;
            STATE_0A5B: if (cnt==11'd45) cnt <= 0; else cnt <= cnt + 1;
            STATE_0A3B: if (cnt==11'd1921) cnt <= 0; else cnt <= cnt + 1;
            STATE_0A2B: if (cnt==11'd781) cnt <= 0; else cnt <= cnt + 1;
            STATE_OUTPUT: if (cnt==11'd4) cnt <= 0; else cnt <= cnt + 1;
            default: cnt <= 11'd0;
        endcase
end

// Store Input
always @(posedge clk or negedge rst_n) begin // read 1st keyboard
    if (!rst_n) keyboard_arr[0] <= 0;
    else
    case (current_state)
        STATE_IDLE: if (in_valid) keyboard_arr[0] <= keyboard; else keyboard_arr[0] <= keyboard_arr[0];
        default: keyboard_arr[0] <= keyboard_arr[0];
    endcase
end

generate // read 2-8th keyboard
    for (vi=1;vi<8;vi=vi+1) begin: keyboard_2_to_7
        always @(posedge clk or negedge rst_n) begin 
            if (!rst_n) keyboard_arr[vi] <= 0;
            else
            case (current_state)
                STATE_INPUT: if (cnt==vi-1) keyboard_arr[vi] <= keyboard; else keyboard_arr[vi] <= keyboard_arr[vi];
                default: keyboard_arr[vi] <= keyboard_arr[vi];
            endcase
        end
    end
endgenerate

always @(posedge clk or negedge rst_n) begin // read 1st answer
    if (!rst_n) begin
        answer_arr[0] <= 0;
    end
    else
    case (current_state)
        STATE_IDLE: if (in_valid) answer_arr[0] <= answer; else answer_arr[0] <= answer_arr[0];
        default: answer_arr[0] <= answer_arr[0];
    endcase
end

always @(posedge clk or negedge rst_n) begin // read 2nd answer
    if (!rst_n) begin
        answer_arr[1] <= 0;
    end
    else
    case (current_state)
        STATE_INPUT: if (cnt==0) answer_arr[1] <= answer; else answer_arr[1] <= answer_arr[1]; 
        default: answer_arr[1] <= answer_arr[1];
    endcase
end

always @(posedge clk or negedge rst_n) begin // read 3rd answer
    if (!rst_n) begin
        answer_arr[2] <= 0;
    end
    else
    case (current_state)
        STATE_INPUT: if (cnt==1) answer_arr[2] <= answer; else answer_arr[2] <= answer_arr[2]; 
        default: answer_arr[2] <= answer_arr[2];
    endcase
end

always @(posedge clk or negedge rst_n) begin // read 4th answer
    if (!rst_n) begin
        answer_arr[3] <= 0;
    end
    else
    case (current_state)
        STATE_INPUT: if (cnt==2) answer_arr[3] <= answer; else answer_arr[3] <= answer_arr[3]; 
        default: answer_arr[3] <= answer_arr[3];
    endcase
end

always @(posedge clk or negedge rst_n) begin // read 5th answer
    if (!rst_n) begin
        answer_arr[4] <= 0;
    end
    else
    case (current_state)
        STATE_INPUT: if (cnt==3) answer_arr[4] <= answer; else answer_arr[4] <= answer_arr[4]; 
        default: answer_arr[4] <= answer_arr[4];
    endcase
end

// generate // read 2-5th answer
//     for (vi=1;vi<5;vi=vi+1) begin: answer_2_to_4
//         always @(posedge clk or negedge rst_n) begin
//             if (!rst_n) answer_arr[vi] <= 0;
//             else
//             case (current_state)
//                 STATE_INPUT: if (cnt==vi-1) answer_arr[vi] <= answer; else answer_arr[vi] <= answer[vi];
//                 default: answer_arr[vi] <= answer_arr[vi];
//             endcase
//         end
//     end
// endgenerate

always @(posedge clk or negedge rst_n) begin // read 1st weight
    if (!rst_n) begin
        weight_arr[0] <= 0;
    end
    else
    case (current_state)
        STATE_IDLE: if (in_valid) weight_arr[0] <= weight; else weight_arr[0] <= weight_arr[0];
        default: weight_arr[0] <= weight_arr[0];
    endcase
end

generate // read 2-5th weight
    for (vi=1;vi<5;vi=vi+1) begin: weight_2_to_4
        always @(posedge clk or negedge rst_n) begin
            if (!rst_n) weight_arr[vi] <= 0;
            else
            case (current_state)
                STATE_INPUT: if (cnt==vi-1) weight_arr[vi] <= weight; else weight_arr[vi] <= weight_arr[vi];
                default: weight_arr[vi] <= weight_arr[vi];
            endcase
        end
    end
endgenerate

always @(posedge clk or negedge rst_n) begin // read 1st match_target
    if (!rst_n) begin
        match_target_arr[0] <= 0;
    end
    else
    case (current_state)
        STATE_IDLE: if (in_valid) match_target_arr[0] <= match_target; else match_target_arr[0] <= match_target_arr[0];
        default: match_target_arr[0] <= match_target_arr[0];
    endcase
end

always @(posedge clk or negedge rst_n) begin // read 2nd match_target
    if (!rst_n) begin
        match_target_arr[1] <= 0;
    end
    else
    case (current_state)
        STATE_INPUT: if (cnt==0) match_target_arr[1] <= match_target; else match_target_arr[1] <= match_target_arr[1];
        default: match_target_arr[1] <= match_target_arr[1];
    endcase
end

always @(posedge clk or negedge rst_n) begin // reorder sequence along answer sequence (resource sharing TBD)
    if (!rst_n) begin
        for (ii=0;ii<8;ii=ii+1) begin
            reorder_arr[ii] <= 0;
        end
    end
    else case (current_state)
        STATE_REORDER:
            case (cnt)
                0: begin
                    reorder_arr[0] <= keyboard_arr[0]; 
                    reorder_arr[1] <= keyboard_arr[1]; 
                    reorder_arr[2] <= keyboard_arr[2]; 
                    reorder_arr[3] <= keyboard_arr[3]; 
                    reorder_arr[4] <= keyboard_arr[4]; 
                    reorder_arr[5] <= keyboard_arr[5]; 
                    reorder_arr[6] <= keyboard_arr[6];
                    reorder_arr[7] <= keyboard_arr[7];           
                end
                1: if (answer_arr[0]==reorder_arr[1]) begin reorder_arr[0] <= reorder_arr[1]; reorder_arr[1] <= reorder_arr[0]; end
                2: if (answer_arr[0]==reorder_arr[2]) begin reorder_arr[0] <= reorder_arr[2]; reorder_arr[2] <= reorder_arr[0]; end
                3: if (answer_arr[0]==reorder_arr[3]) begin reorder_arr[0] <= reorder_arr[3]; reorder_arr[3] <= reorder_arr[0]; end
                4: if (answer_arr[0]==reorder_arr[4]) begin reorder_arr[0] <= reorder_arr[4]; reorder_arr[4] <= reorder_arr[0]; end
                5: if (answer_arr[0]==reorder_arr[5]) begin reorder_arr[0] <= reorder_arr[5]; reorder_arr[5] <= reorder_arr[0]; end
                6: if (answer_arr[0]==reorder_arr[6]) begin reorder_arr[0] <= reorder_arr[6]; reorder_arr[6] <= reorder_arr[0]; end
                7: if (answer_arr[0]==reorder_arr[7]) begin reorder_arr[0] <= reorder_arr[7]; reorder_arr[7] <= reorder_arr[0]; end

                8: if (answer_arr[1]==reorder_arr[2]) begin reorder_arr[1] <= reorder_arr[2]; reorder_arr[2] <= reorder_arr[1]; end
                9: if (answer_arr[1]==reorder_arr[3]) begin reorder_arr[1] <= reorder_arr[3]; reorder_arr[3] <= reorder_arr[1]; end
                10: if (answer_arr[1]==reorder_arr[4]) begin reorder_arr[1] <= reorder_arr[4]; reorder_arr[4] <= reorder_arr[1]; end
                11: if (answer_arr[1]==reorder_arr[5]) begin reorder_arr[1] <= reorder_arr[5]; reorder_arr[5] <= reorder_arr[1]; end
                12: if (answer_arr[1]==reorder_arr[6]) begin reorder_arr[1] <= reorder_arr[6]; reorder_arr[6] <= reorder_arr[1]; end
                13: if (answer_arr[1]==reorder_arr[7]) begin reorder_arr[1] <= reorder_arr[7]; reorder_arr[7] <= reorder_arr[1]; end

                14: if (answer_arr[2]==reorder_arr[3]) begin reorder_arr[2] <= reorder_arr[3]; reorder_arr[3] <= reorder_arr[2]; end
                15: if (answer_arr[2]==reorder_arr[4]) begin reorder_arr[2] <= reorder_arr[4]; reorder_arr[4] <= reorder_arr[2]; end
                16: if (answer_arr[2]==reorder_arr[5]) begin reorder_arr[2] <= reorder_arr[5]; reorder_arr[5] <= reorder_arr[2]; end
                17: if (answer_arr[2]==reorder_arr[6]) begin reorder_arr[2] <= reorder_arr[6]; reorder_arr[6] <= reorder_arr[2]; end
                18: if (answer_arr[2]==reorder_arr[7]) begin reorder_arr[2] <= reorder_arr[7]; reorder_arr[7] <= reorder_arr[2]; end

                19: if (answer_arr[3]==reorder_arr[4]) begin reorder_arr[3] <= reorder_arr[4]; reorder_arr[4] <= reorder_arr[3]; end
                20: if (answer_arr[3]==reorder_arr[5]) begin reorder_arr[3] <= reorder_arr[5]; reorder_arr[5] <= reorder_arr[3]; end
                21: if (answer_arr[3]==reorder_arr[6]) begin reorder_arr[3] <= reorder_arr[6]; reorder_arr[6] <= reorder_arr[3]; end
                22: if (answer_arr[3]==reorder_arr[7]) begin reorder_arr[3] <= reorder_arr[7]; reorder_arr[7] <= reorder_arr[3]; end

                23: if (answer_arr[4]==reorder_arr[5]) begin reorder_arr[4] <= reorder_arr[5]; reorder_arr[5] <= reorder_arr[4]; end
                24: if (answer_arr[4]==reorder_arr[6]) begin reorder_arr[4] <= reorder_arr[6]; reorder_arr[6] <= reorder_arr[4]; end
                25: if (answer_arr[4]==reorder_arr[7]) begin reorder_arr[4] <= reorder_arr[7]; reorder_arr[7] <= reorder_arr[4]; end
                default: begin
                    reorder_arr[0] <= reorder_arr[0];
                    reorder_arr[1] <= reorder_arr[1];
                    reorder_arr[2] <= reorder_arr[2];
                    reorder_arr[3] <= reorder_arr[3];
                    reorder_arr[4] <= reorder_arr[4];
                    reorder_arr[5] <= reorder_arr[5];
                    reorder_arr[6] <= reorder_arr[6];
                    reorder_arr[7] <= reorder_arr[7];
                end
            endcase
        default: begin
            reorder_arr[0] <= reorder_arr[0];
            reorder_arr[1] <= reorder_arr[1];
            reorder_arr[2] <= reorder_arr[2];
            reorder_arr[3] <= reorder_arr[3];
            reorder_arr[4] <= reorder_arr[4];
            reorder_arr[5] <= reorder_arr[5];
            reorder_arr[6] <= reorder_arr[6];
            reorder_arr[7] <= reorder_arr[7];
        end
    endcase

end

always @(posedge clk or negedge rst_n) begin // iterating all permutations according to NANB
    if (!rst_n) begin
        // for (ii=0;ii<5;ii=ii+1) begin
        //     perm_arr[ii] <= 0;
        // end
        perm_arr[0] <= 0;
        perm_arr[1] <= 0;
        perm_arr[2] <= 0;
        perm_arr[3] <= 0;
        perm_arr[4] <= 0;
    end
    else
    case (current_state)
        STATE_5A0B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_4A0B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            2: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            3: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            4: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            5: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            7: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            8: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            9: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            10: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            11: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            12: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            13: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            14: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_3A2B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            2: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            3: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            4: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            5: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            7: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            8: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            9: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_3A1B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            2: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            3: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            4: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            5: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            7: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            8: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            9: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            10: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            11: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            12: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            13: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            14: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            15: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            16: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            17: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            18: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            19: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            20: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            21: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            22: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            23: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            24: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            25: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            26: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            27: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            28: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            29: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            30: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            31: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            32: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            33: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            34: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            35: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            36: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            37: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            38: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            39: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            40: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            41: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            42: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            43: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            44: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            45: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            46: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            47: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            48: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            49: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            50: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            51: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            52: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            53: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            54: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            55: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            56: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            57: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            58: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            59: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_3A0B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            2: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            3: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            4: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            5: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            7: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            8: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            9: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            10: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            11: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            12: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            13: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            14: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            15: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            16: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            17: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            18: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            19: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            20: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            21: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            22: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            23: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            24: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            25: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            26: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            27: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            28: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            29: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            30: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            31: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            32: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            33: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            34: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            35: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            36: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            37: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            38: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            39: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            40: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            41: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            42: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            43: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            44: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            45: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            46: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            47: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            48: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            49: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            50: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            51: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            52: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            53: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            54: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            55: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            56: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            57: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            58: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            59: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_2A2B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            1: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            2: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            3: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            4: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            5: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            7: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            8: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            9: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            10: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            11: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            12: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            13: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            14: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            15: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            16: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            17: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            18: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            19: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            20: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            21: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            22: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            23: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            24: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            25: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            26: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            27: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            28: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            29: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            30: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            31: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            32: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            33: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            34: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            35: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            36: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            37: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            38: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            39: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            40: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            41: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            42: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            43: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            44: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            45: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            46: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            47: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            48: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            49: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            50: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            51: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            52: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            53: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            54: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            55: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            56: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            57: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            58: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            59: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            60: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            61: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            62: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            63: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            64: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            65: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            66: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            67: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            68: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            69: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            70: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            71: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            72: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            73: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            74: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            75: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            76: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            77: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            78: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            79: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            80: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            81: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            82: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            83: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            84: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            85: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            86: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            87: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            88: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            89: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            90: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            91: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            92: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            93: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            94: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            95: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            96: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            97: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            98: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            99: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            100: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            101: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            102: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            103: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            104: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            105: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            106: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            107: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            108: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            109: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            110: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            111: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            112: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            113: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            114: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            115: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            116: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            117: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            118: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            119: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            120: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            121: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            122: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            123: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            124: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            125: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            126: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            127: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            128: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            129: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            130: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            131: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            132: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            133: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            134: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            135: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            136: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            137: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            138: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            139: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            140: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            141: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            142: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            143: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            144: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            145: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            146: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            147: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            148: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            149: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            150: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            151: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            152: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            153: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            154: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            155: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            156: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            157: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            158: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            159: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            160: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            161: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            162: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            163: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            164: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            165: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            166: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            167: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            168: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            169: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            170: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            171: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            172: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            173: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            174: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            175: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            176: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            177: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            178: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            179: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            180: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            181: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            182: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            183: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            184: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            185: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            186: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            187: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            188: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            189: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            190: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            191: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            192: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            193: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            194: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            195: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            196: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            197: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            198: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            199: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            200: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            201: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            202: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            203: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            204: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            205: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            206: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            207: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            208: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            209: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            210: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            211: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            212: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            213: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            214: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            215: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            216: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            217: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            218: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            219: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            220: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            221: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            222: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            223: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            224: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            225: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            226: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            227: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            228: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            229: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            230: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            231: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            232: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            233: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            234: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            235: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            236: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            237: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            238: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            239: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            240: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            241: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            242: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            243: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            244: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            245: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            246: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            247: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            248: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            249: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            250: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            251: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            252: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            253: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            254: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            255: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            256: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            257: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            258: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            259: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            260: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            261: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            262: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            263: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            264: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            265: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            266: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            267: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            268: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            269: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_2A3B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            2: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            3: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            4: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            5: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            7: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            8: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            9: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            10: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            11: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            12: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            13: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            14: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            15: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            16: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            17: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            18: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            19: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_2A1B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            1: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            2: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            3: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            4: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            5: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            7: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            8: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            9: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            10: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            11: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            12: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            13: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            14: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            15: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            16: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            17: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            18: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            19: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            20: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            21: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            22: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            23: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            24: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            25: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            26: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            27: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            28: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            29: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            30: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            31: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            32: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            33: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            34: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            35: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            36: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            37: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            38: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            39: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            40: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            41: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            42: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            43: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            44: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            45: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            46: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            47: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            48: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            49: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            50: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            51: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            52: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            53: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            54: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            55: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            56: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            57: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            58: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            59: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            60: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            61: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            62: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            63: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            64: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            65: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            66: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            67: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            68: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            69: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            70: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            71: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            72: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            73: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            74: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            75: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            76: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            77: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            78: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            79: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            80: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            81: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            82: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            83: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            84: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            85: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            86: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            87: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            88: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            89: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            90: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            91: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            92: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            93: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            94: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            95: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            96: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            97: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            98: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            99: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            100: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            101: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            102: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            103: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            104: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            105: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            106: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            107: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            108: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            109: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            110: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            111: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            112: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            113: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            114: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            115: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            116: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            117: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            118: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            119: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            120: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            121: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            122: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            123: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            124: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            125: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            126: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            127: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            128: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            129: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            130: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            131: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            132: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            133: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            134: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            135: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            136: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            137: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            138: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            139: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            140: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            141: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            142: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            143: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            144: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            145: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            146: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            147: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            148: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            149: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            150: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            151: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            152: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            153: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            154: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            155: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            156: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            157: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            158: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            159: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            160: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            161: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            162: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            163: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            164: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            165: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            166: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            167: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            168: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            169: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            170: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            171: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            172: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            173: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            174: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            175: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            176: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            177: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            178: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            179: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            180: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            181: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            182: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            183: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            184: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            185: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            186: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            187: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            188: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            189: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            190: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            191: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            192: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            193: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            194: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            195: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            196: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            197: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            198: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            199: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            200: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            201: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            202: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            203: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            204: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            205: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            206: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            207: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            208: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            209: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            210: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            211: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            212: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            213: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            214: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            215: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            216: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            217: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            218: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            219: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            220: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            221: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            222: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            223: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            224: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            225: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            226: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            227: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            228: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            229: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            230: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            231: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            232: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            233: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            234: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            235: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            236: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            237: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            238: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            239: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            240: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            241: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            242: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            243: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            244: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            245: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            246: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            247: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            248: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            249: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            250: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            251: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            252: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            253: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            254: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            255: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            256: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            257: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            258: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            259: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            260: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            261: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            262: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            263: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            264: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            265: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            266: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            267: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            268: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            269: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            270: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            271: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            272: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            273: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            274: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            275: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            276: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            277: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            278: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            279: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            280: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            281: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            282: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            283: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            284: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            285: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            286: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            287: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            288: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            289: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            290: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            291: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            292: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            293: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            294: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            295: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            296: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            297: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            298: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            299: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            300: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            301: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            302: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            303: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            304: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            305: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            306: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            307: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            308: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            309: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            310: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            311: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            312: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            313: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            314: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            315: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            316: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            317: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            318: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            319: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            320: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            321: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            322: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            323: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            324: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            325: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            326: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            327: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            328: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            329: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            330: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            331: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            332: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            333: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            334: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            335: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            336: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            337: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            338: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            339: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            340: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            341: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            342: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            343: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            344: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            345: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            346: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            347: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            348: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            349: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            350: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            351: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            352: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            353: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            354: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            355: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            356: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            357: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            358: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            359: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_2A0B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            1: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            2: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            3: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            4: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            5: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            6: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            7: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            8: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            9: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            10: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            11: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            12: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            13: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            14: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            15: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            16: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            17: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            18: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            19: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            20: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            21: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            22: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            23: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            24: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            25: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            26: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            27: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            28: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            29: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            30: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            31: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            32: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            33: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            34: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            35: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            36: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            37: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            38: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            39: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            40: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            41: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            42: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            43: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            44: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            45: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            46: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            47: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            48: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            49: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            50: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            51: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            52: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            53: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            54: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            55: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            56: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            57: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[4]; end
            58: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            59: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_1A4B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            2: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            3: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            4: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            5: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            6: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            7: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            8: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            9: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            10: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            11: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            12: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            13: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            14: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            15: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            16: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            17: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            18: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            19: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            20: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            21: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            22: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            23: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            24: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            25: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            26: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            27: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            28: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            29: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            30: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            31: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            32: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            33: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            34: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            35: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            36: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            37: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            38: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            39: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            40: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            41: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            42: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            43: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            44: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_1A3B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            2: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            3: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            4: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            5: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            6: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            7: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            8: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            9: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            10: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            11: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            12: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            13: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            14: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            15: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            16: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            17: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            18: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            19: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            20: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            21: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            22: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            23: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            24: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            25: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            26: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            27: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            28: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            29: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            30: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            31: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            32: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            33: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            34: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            35: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            36: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            37: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            38: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            39: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            40: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            41: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            42: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            43: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            44: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            45: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            46: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            47: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            48: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            49: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            50: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            51: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            52: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            53: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            54: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            55: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            56: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            57: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            58: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            59: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            60: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            61: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            62: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            63: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            64: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            65: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            66: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            67: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            68: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            69: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            70: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            71: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            72: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            73: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            74: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            75: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            76: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            77: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            78: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            79: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            80: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            81: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            82: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            83: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            84: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            85: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            86: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            87: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            88: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            89: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            90: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            91: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            92: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            93: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            94: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            95: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            96: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            97: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            98: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            99: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            100: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            101: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            102: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            103: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            104: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            105: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            106: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            107: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            108: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            109: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            110: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            111: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            112: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            113: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            114: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            115: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            116: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            117: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            118: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            119: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            120: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            121: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            122: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            123: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            124: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            125: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            126: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            127: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            128: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            129: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            130: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            131: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            132: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            133: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            134: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            135: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            136: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            137: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            138: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            139: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            140: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            141: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            142: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            143: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            144: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            145: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            146: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            147: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            148: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            149: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            150: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            151: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            152: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            153: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            154: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            155: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            156: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            157: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            158: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            159: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            160: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            161: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            162: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            163: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            164: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            165: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            166: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            167: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            168: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            169: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            170: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            171: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            172: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            173: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            174: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            175: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            176: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            177: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            178: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            179: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            180: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            181: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            182: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            183: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            184: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            185: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            186: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            187: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            188: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            189: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            190: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            191: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            192: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            193: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            194: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            195: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            196: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            197: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            198: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            199: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            200: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            201: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            202: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            203: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            204: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            205: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            206: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            207: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            208: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            209: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            210: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            211: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            212: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            213: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            214: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            215: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            216: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            217: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            218: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            219: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            220: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            221: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            222: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            223: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            224: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            225: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            226: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            227: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            228: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            229: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            230: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            231: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            232: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            233: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            234: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            235: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            236: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            237: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            238: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            239: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            240: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            241: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            242: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            243: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            244: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            245: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            246: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            247: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            248: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            249: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            250: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            251: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            252: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            253: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            254: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            255: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            256: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            257: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            258: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            259: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            260: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            261: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            262: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            263: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            264: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            265: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            266: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            267: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            268: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            269: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            270: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            271: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            272: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            273: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            274: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            275: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            276: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            277: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            278: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            279: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            280: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            281: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            282: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            283: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            284: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            285: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            286: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            287: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            288: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            289: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            290: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            291: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            292: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            293: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            294: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            295: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            296: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            297: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            298: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            299: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            300: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            301: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            302: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            303: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            304: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            305: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            306: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            307: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            308: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            309: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            310: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            311: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            312: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            313: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            314: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            315: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            316: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            317: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            318: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            319: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            320: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            321: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            322: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            323: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            324: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            325: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            326: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            327: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            328: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            329: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            330: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            331: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            332: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            333: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            334: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            335: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            336: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            337: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            338: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            339: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            340: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            341: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            342: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            343: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            344: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            345: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            346: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            347: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            348: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            349: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            350: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            351: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            352: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            353: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            354: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            355: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            356: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            357: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            358: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            359: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            360: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            361: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            362: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            363: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            364: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            365: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            366: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            367: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            368: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            369: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            370: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            371: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            372: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            373: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            374: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            375: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            376: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            377: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            378: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            379: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            380: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            381: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            382: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            383: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            384: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            385: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            386: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            387: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            388: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            389: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            390: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            391: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            392: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            393: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            394: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            395: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            396: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            397: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            398: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            399: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            400: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            401: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            402: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            403: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            404: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            405: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            406: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            407: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            408: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            409: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            410: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            411: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            412: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            413: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            414: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            415: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            416: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            417: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            418: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            419: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            420: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            421: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            422: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            423: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            424: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            425: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            426: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            427: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            428: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            429: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            430: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            431: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            432: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            433: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            434: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            435: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            436: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            437: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            438: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            439: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            440: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            441: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            442: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            443: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            444: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            445: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            446: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            447: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            448: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            449: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            450: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            451: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            452: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            453: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            454: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            455: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            456: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            457: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            458: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            459: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            460: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            461: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            462: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            463: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            464: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            465: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            466: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            467: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            468: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            469: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            470: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            471: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            472: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            473: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            474: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            475: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            476: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            477: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            478: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            479: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            480: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            481: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            482: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            483: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            484: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            485: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            486: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            487: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            488: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            489: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            490: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            491: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            492: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            493: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            494: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            495: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            496: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            497: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            498: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            499: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            500: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            501: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            502: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            503: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            504: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            505: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            506: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            507: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            508: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            509: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            510: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            511: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            512: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            513: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            514: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            515: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            516: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            517: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            518: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            519: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            520: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            521: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            522: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            523: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            524: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            525: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            526: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            527: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            528: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            529: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            530: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            531: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            532: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            533: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            534: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            535: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            536: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            537: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            538: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            539: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            540: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            541: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            542: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            543: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            544: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            545: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            546: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            547: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            548: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            549: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            550: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            551: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            552: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            553: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            554: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            555: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            556: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            557: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            558: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            559: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            560: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            561: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            562: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            563: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            564: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            565: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            566: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            567: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            568: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            569: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            570: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            571: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            572: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            573: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            574: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            575: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            576: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            577: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            578: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            579: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            580: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            581: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            582: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            583: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            584: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            585: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            586: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            587: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            588: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            589: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            590: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            591: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            592: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            593: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            594: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            595: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            596: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            597: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            598: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            599: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            600: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            601: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            602: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            603: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            604: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            605: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            606: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            607: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            608: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            609: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            610: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            611: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            612: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            613: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            614: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            615: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            616: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            617: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            618: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            619: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            620: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            621: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            622: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            623: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            624: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            625: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            626: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            627: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            628: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            629: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            630: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            631: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            632: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            633: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            634: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            635: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            636: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            637: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            638: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            639: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            640: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            641: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            642: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            643: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            644: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            645: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            646: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            647: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            648: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            649: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            650: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            651: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            652: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            653: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            654: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            655: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            656: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            657: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            658: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            659: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_1A2B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            1: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            2: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            3: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            4: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            5: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            6: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            7: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            8: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            9: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            10: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            11: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            12: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            13: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            14: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            15: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            16: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            17: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            18: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            19: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            20: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            21: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            22: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            23: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            24: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            25: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            26: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            27: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            28: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            29: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            30: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            31: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            32: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            33: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            34: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            35: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            36: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            37: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            38: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            39: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            40: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            41: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            42: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            43: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            44: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            45: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            46: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            47: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            48: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            49: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            50: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            51: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            52: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            53: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            54: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            55: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            56: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            57: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            58: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            59: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            60: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            61: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            62: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            63: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            64: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            65: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            66: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            67: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            68: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            69: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            70: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            71: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            72: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            73: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            74: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            75: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            76: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            77: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            78: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            79: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            80: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            81: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            82: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            83: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            84: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            85: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            86: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            87: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            88: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            89: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            90: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            91: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            92: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            93: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            94: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            95: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            96: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            97: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            98: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            99: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            100: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            101: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            102: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            103: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            104: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            105: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            106: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            107: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            108: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            109: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            110: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            111: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            112: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            113: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            114: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            115: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            116: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            117: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            118: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            119: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            120: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            121: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            122: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            123: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            124: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            125: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            126: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            127: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            128: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            129: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            130: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            131: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            132: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            133: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            134: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            135: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            136: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            137: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            138: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            139: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            140: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            141: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            142: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            143: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            144: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            145: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            146: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            147: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            148: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            149: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            150: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            151: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            152: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            153: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            154: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            155: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            156: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            157: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            158: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            159: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            160: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            161: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            162: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            163: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            164: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            165: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            166: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            167: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            168: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            169: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            170: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            171: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            172: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            173: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            174: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            175: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            176: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            177: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            178: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            179: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            180: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            181: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            182: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            183: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            184: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            185: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            186: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            187: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            188: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            189: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            190: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            191: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            192: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            193: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            194: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            195: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            196: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            197: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            198: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            199: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            200: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            201: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            202: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            203: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            204: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            205: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            206: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            207: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            208: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            209: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            210: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            211: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            212: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            213: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            214: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            215: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            216: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            217: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            218: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            219: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            220: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            221: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            222: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            223: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            224: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            225: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            226: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            227: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            228: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            229: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            230: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            231: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            232: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            233: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            234: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            235: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            236: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            237: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            238: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            239: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            240: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            241: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            242: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            243: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            244: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            245: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            246: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            247: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            248: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            249: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            250: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            251: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            252: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            253: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            254: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            255: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            256: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            257: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            258: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            259: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            260: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            261: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            262: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            263: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            264: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            265: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            266: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            267: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            268: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            269: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            270: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            271: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            272: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            273: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            274: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            275: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            276: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            277: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            278: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            279: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            280: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            281: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            282: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            283: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            284: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            285: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            286: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            287: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            288: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            289: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            290: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            291: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            292: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            293: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            294: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            295: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            296: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            297: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            298: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            299: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            300: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            301: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            302: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            303: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            304: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            305: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            306: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            307: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            308: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            309: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            310: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            311: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            312: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            313: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            314: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            315: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            316: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            317: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            318: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            319: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            320: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            321: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            322: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            323: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            324: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            325: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            326: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            327: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            328: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            329: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            330: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            331: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            332: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            333: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            334: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            335: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            336: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            337: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            338: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            339: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            340: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            341: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            342: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            343: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            344: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            345: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            346: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            347: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            348: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            349: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            350: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            351: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            352: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            353: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            354: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            355: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            356: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            357: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            358: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            359: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            360: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            361: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            362: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            363: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            364: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            365: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            366: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            367: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            368: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            369: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            370: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            371: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            372: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            373: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            374: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            375: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            376: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            377: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            378: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            379: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            380: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            381: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            382: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            383: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            384: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            385: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            386: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            387: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            388: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            389: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            390: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            391: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            392: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            393: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            394: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            395: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            396: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            397: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            398: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            399: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            400: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            401: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            402: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            403: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            404: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            405: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            406: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            407: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            408: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            409: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            410: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            411: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            412: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            413: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            414: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            415: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            416: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            417: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            418: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            419: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            420: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            421: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            422: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            423: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            424: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            425: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            426: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            427: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            428: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            429: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            430: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            431: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            432: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            433: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            434: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            435: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            436: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            437: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            438: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            439: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            440: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            441: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            442: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            443: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            444: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            445: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            446: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            447: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            448: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            449: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            450: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            451: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            452: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            453: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            454: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            455: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            456: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            457: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            458: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            459: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            460: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            461: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            462: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            463: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            464: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            465: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            466: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            467: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            468: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            469: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            470: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            471: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            472: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            473: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            474: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            475: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            476: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            477: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            478: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            479: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            480: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            481: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            482: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            483: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            484: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            485: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            486: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            487: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            488: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            489: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            490: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            491: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            492: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            493: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            494: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            495: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            496: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            497: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            498: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            499: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            500: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            501: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            502: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            503: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            504: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            505: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            506: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            507: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            508: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            509: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            510: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            511: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            512: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            513: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            514: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            515: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            516: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            517: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            518: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            519: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            520: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            521: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            522: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            523: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            524: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            525: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            526: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            527: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            528: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            529: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            530: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            531: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            532: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            533: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            534: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            535: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            536: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            537: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            538: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            539: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            540: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            541: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            542: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            543: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            544: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            545: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            546: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            547: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            548: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            549: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            550: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            551: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            552: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            553: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            554: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            555: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            556: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            557: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            558: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            559: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            560: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            561: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            562: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            563: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            564: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            565: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            566: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            567: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            568: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            569: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            570: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            571: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            572: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            573: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            574: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            575: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            576: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            577: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            578: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            579: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            580: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            581: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            582: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            583: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            584: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            585: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            586: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            587: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            588: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            589: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            590: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            591: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            592: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            593: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            594: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            595: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            596: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            597: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            598: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            599: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            600: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            601: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            602: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            603: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            604: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            605: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            606: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            607: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            608: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            609: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            610: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            611: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            612: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            613: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            614: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            615: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            616: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            617: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            618: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            619: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            620: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            621: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            622: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            623: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            624: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            625: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            626: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            627: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            628: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            629: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            630: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            631: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            632: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            633: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            634: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            635: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            636: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            637: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            638: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            639: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            640: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            641: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            642: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            643: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            644: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            645: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            646: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            647: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            648: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            649: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            650: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            651: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            652: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            653: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            654: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            655: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            656: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            657: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            658: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            659: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            660: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            661: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            662: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            663: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            664: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            665: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            666: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            667: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            668: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            669: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            670: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            671: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            672: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            673: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            674: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            675: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            676: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            677: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            678: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            679: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            680: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            681: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            682: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            683: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            684: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            685: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            686: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            687: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            688: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            689: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            690: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            691: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            692: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            693: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            694: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            695: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            696: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            697: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            698: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            699: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            700: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            701: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            702: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            703: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            704: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            705: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            706: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            707: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            708: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            709: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            710: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            711: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            712: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            713: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            714: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            715: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            716: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            717: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            718: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            719: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            720: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            721: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            722: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            723: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            724: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            725: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            726: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            727: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            728: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            729: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            730: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            731: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            732: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            733: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            734: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            735: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            736: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            737: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            738: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            739: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            740: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            741: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            742: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            743: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            744: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            745: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            746: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            747: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            748: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            749: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            750: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            751: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            752: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            753: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            754: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            755: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            756: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            757: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            758: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            759: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            760: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            761: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            762: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            763: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            764: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            765: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            766: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            767: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            768: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            769: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            770: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            771: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            772: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            773: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            774: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            775: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            776: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            777: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            778: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            779: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            780: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            781: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            782: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            783: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            784: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            785: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            786: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            787: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            788: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            789: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            790: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            791: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            792: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            793: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            794: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            795: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            796: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            797: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            798: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            799: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            800: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            801: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            802: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            803: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            804: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            805: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            806: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            807: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            808: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            809: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            810: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            811: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            812: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            813: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            814: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            815: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            816: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            817: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            818: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            819: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            820: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            821: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            822: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            823: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            824: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            825: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            826: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            827: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            828: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            829: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            830: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            831: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            832: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            833: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            834: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            835: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            836: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            837: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            838: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            839: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            840: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            841: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            842: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            843: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            844: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            845: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            846: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            847: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            848: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            849: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            850: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            851: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            852: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            853: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            854: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            855: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            856: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            857: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            858: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            859: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            860: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            861: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            862: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            863: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            864: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            865: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            866: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            867: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            868: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            869: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            870: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            871: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            872: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            873: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            874: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            875: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            876: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            877: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            878: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            879: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            880: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            881: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            882: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            883: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            884: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            885: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            886: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            887: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            888: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            889: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            890: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            891: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            892: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            893: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            894: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            895: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            896: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            897: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            898: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            899: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            900: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            901: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            902: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            903: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            904: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            905: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            906: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            907: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            908: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            909: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            910: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            911: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            912: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            913: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            914: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            915: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            916: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            917: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            918: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            919: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            920: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            921: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            922: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            923: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            924: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            925: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            926: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            927: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            928: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            929: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            930: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            931: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            932: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            933: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            934: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            935: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            936: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            937: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            938: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            939: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            940: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            941: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            942: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            943: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            944: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            945: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            946: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            947: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            948: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            949: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            950: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            951: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            952: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            953: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            954: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            955: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            956: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            957: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            958: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            959: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            960: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            961: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            962: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            963: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            964: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            965: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            966: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            967: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            968: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            969: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            970: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            971: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            972: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            973: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            974: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            975: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            976: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            977: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            978: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            979: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            980: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            981: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            982: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            983: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            984: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            985: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            986: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            987: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            988: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            989: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            990: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            991: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            992: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            993: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            994: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            995: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            996: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            997: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            998: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            999: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            1000: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1001: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            1002: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1003: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1004: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1005: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1006: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1007: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1008: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1009: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1010: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1011: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            1012: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1013: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            1014: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1015: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1016: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1017: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1018: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1019: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1020: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1021: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1022: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1023: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1024: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1025: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1026: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1027: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1028: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1029: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1030: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1031: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            1032: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1033: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            1034: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1035: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1036: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1037: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1038: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1039: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1040: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1041: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1042: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1043: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1044: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1045: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1046: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1047: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1048: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1049: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1050: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1051: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1052: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1053: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1054: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1055: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1056: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1057: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1058: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1059: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1060: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1061: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1062: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1063: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1064: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1065: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1066: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1067: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1068: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1069: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1070: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1071: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1072: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1073: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1074: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1075: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1076: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1077: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1078: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1079: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1080: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1081: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1082: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1083: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1084: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1085: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1086: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1087: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1088: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1089: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1090: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1091: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1092: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1093: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            1094: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1095: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1096: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1097: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1098: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1099: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1100: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1101: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1102: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1103: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1104: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1105: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1106: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1107: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            1108: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1109: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1110: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1111: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1112: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1113: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1114: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1115: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1116: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1117: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1118: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1119: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1120: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1121: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1122: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1123: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1124: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1125: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1126: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1127: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1128: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1129: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1130: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1131: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1132: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1133: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1134: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1135: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1136: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1137: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1138: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1139: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1140: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1141: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1142: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1143: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1144: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1145: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1146: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1147: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1148: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1149: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1150: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1151: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1152: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1153: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1154: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1155: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1156: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1157: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1158: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1159: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            1160: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1161: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1162: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1163: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            1164: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1165: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1166: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1167: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1168: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1169: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            1170: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1171: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1172: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1173: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1174: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1175: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1176: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1177: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1178: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1179: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1180: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            1181: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            1182: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1183: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1184: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1185: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1186: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1187: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1188: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1189: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1190: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1191: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1192: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1193: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1194: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1195: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1196: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1197: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1198: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1199: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            1200: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            1201: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            1202: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1203: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1204: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1205: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1206: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1207: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1208: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1209: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1210: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1211: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1212: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1213: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1214: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1215: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1216: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1217: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1218: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1219: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1220: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1221: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1222: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1223: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1224: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1225: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1226: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1227: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1228: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1229: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1230: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1231: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1232: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1233: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1234: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1235: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1236: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1237: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1238: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1239: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1240: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1241: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1242: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1243: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1244: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1245: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1246: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            1247: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1248: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1249: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1250: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1251: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1252: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1253: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1254: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            1255: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            1256: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            1257: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            1258: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            1259: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_1A1B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            1: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            2: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            3: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            4: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            5: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            6: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            7: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            8: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            9: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            10: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            11: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            12: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            13: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            14: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            15: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            16: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            17: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            18: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            19: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            20: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            21: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            22: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            23: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            24: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            25: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            26: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            27: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            28: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            29: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            30: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            31: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            32: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            33: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            34: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            35: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            36: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            37: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            38: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            39: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            40: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            41: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            42: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            43: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            44: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            45: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            46: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            47: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            48: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            49: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            50: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            51: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            52: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            53: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            54: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            55: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            56: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            57: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            58: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            59: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            60: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            61: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            62: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            63: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            64: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            65: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            66: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            67: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            68: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            69: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            70: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            71: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            72: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            73: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            74: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            75: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            76: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            77: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            78: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            79: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            80: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            81: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            82: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            83: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            84: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            85: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            86: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            87: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            88: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            89: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            90: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            91: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            92: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            93: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            94: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            95: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            96: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            97: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            98: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            99: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            100: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            101: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            102: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            103: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            104: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            105: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            106: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            107: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            108: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            109: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            110: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            111: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            112: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            113: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            114: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            115: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            116: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            117: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            118: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            119: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            120: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            121: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            122: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            123: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            124: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            125: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            126: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            127: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            128: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            129: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            130: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            131: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            132: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            133: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            134: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            135: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            136: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            137: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            138: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            139: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            140: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            141: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            142: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            143: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            144: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            145: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            146: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            147: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            148: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            149: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            150: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            151: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            152: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            153: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            154: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            155: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            156: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            157: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            158: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            159: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            160: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            161: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            162: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            163: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            164: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            165: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            166: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            167: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            168: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            169: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            170: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            171: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            172: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            173: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            174: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            175: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            176: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            177: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            178: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            179: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            180: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            181: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            182: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            183: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            184: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            185: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            186: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            187: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            188: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            189: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            190: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            191: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            192: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            193: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            194: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            195: begin perm_arr[0]<=reorder_arr[0];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            196: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            197: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            198: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            199: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            200: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            201: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            202: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            203: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            204: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            205: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            206: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            207: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            208: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            209: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            210: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            211: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            212: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            213: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            214: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            215: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            216: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            217: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            218: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            219: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            220: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            221: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            222: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            223: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            224: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            225: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            226: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            227: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            228: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            229: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            230: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            231: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            232: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            233: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            234: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            235: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            236: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            237: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            238: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            239: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            240: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            241: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            242: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            243: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            244: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            245: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            246: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            247: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            248: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            249: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            250: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            251: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            252: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            253: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            254: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            255: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            256: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            257: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            258: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            259: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            260: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            261: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            262: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            263: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            264: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            265: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            266: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            267: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            268: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            269: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            270: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            271: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            272: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            273: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            274: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            275: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            276: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            277: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            278: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            279: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            280: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            281: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            282: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            283: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            284: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            285: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            286: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            287: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            288: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            289: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            290: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            291: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            292: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[4]; end
            293: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            294: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            295: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            296: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            297: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            298: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            299: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            300: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            301: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            302: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            303: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            304: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            305: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            306: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            307: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            308: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            309: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            310: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            311: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            312: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            313: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            314: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            315: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            316: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[4]; end
            317: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[4]; end
            318: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[4]; end
            319: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[0]; end
            320: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[1]; end
            321: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[2]; end
            322: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            323: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            324: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            325: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            326: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            327: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            328: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            329: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[4]; end
            330: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            331: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            332: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            333: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            334: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[4]; end
            335: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[6]; end
            336: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            337: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            338: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            339: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            340: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            341: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            342: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            343: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[2];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            344: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            345: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            346: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            347: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            348: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            349: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            350: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            351: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            352: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[7]; end
            353: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            354: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            355: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            356: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            357: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            358: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[1];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            359: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[3];perm_arr[4]<=reorder_arr[5]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_0A4B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            2: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            3: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            4: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            5: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            6: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            7: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            8: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            9: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            10: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            11: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            12: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            13: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            14: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            15: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            16: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            17: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            18: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            19: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            20: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            21: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            22: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            23: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            24: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            25: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            26: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            27: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            28: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            29: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            30: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            31: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            32: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            33: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            34: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            35: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            36: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            37: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            38: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            39: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            40: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            41: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            42: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            43: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            44: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            45: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            46: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            47: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            48: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            49: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            50: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            51: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            52: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            53: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            54: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            55: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            56: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            57: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            58: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            59: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            60: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            61: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            62: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            63: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            64: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            65: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            66: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            67: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            68: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            69: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            70: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            71: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            72: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            73: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            74: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            75: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            76: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            77: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            78: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            79: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            80: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            81: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            82: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            83: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            84: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            85: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            86: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            87: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            88: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            89: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            90: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            91: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            92: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            93: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            94: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            95: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            96: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            97: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            98: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            99: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            100: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            101: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            102: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            103: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            104: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            105: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            106: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            107: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            108: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            109: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            110: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            111: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            112: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            113: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            114: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            115: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            116: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            117: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            118: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            119: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            120: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            121: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            122: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            123: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            124: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            125: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            126: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            127: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            128: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            129: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            130: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            131: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            132: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            133: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            134: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            135: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            136: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            137: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            138: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            139: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            140: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            141: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            142: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            143: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            144: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            145: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            146: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            147: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            148: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            149: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            150: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            151: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            152: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            153: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            154: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            155: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            156: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            157: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            158: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            159: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            160: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            161: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            162: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            163: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            164: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            165: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            166: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            167: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            168: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            169: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            170: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            171: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            172: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            173: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            174: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            175: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            176: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            177: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            178: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            179: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            180: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            181: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            182: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            183: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            184: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            185: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            186: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            187: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            188: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            189: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            190: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            191: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            192: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            193: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            194: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            195: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            196: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            197: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            198: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            199: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            200: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            201: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            202: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            203: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            204: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            205: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            206: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            207: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            208: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            209: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            210: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            211: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            212: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            213: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            214: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            215: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            216: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            217: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            218: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            219: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            220: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            221: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            222: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            223: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            224: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            225: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            226: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            227: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            228: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            229: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            230: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            231: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            232: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            233: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            234: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            235: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            236: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            237: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            238: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            239: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            240: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            241: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            242: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            243: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            244: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            245: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            246: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            247: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            248: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            249: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            250: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            251: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            252: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            253: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            254: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            255: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            256: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            257: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            258: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            259: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            260: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            261: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            262: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            263: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            264: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            265: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            266: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            267: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            268: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            269: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            270: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            271: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            272: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            273: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            274: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            275: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            276: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            277: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            278: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            279: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            280: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            281: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            282: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            283: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            284: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            285: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            286: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            287: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            288: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            289: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            290: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            291: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            292: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            293: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            294: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            295: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            296: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            297: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            298: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            299: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            300: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            301: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            302: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            303: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            304: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            305: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            306: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            307: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            308: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            309: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            310: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            311: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            312: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            313: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            314: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            315: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            316: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            317: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            318: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            319: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            320: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            321: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            322: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            323: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            324: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            325: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            326: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            327: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            328: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            329: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            330: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            331: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            332: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            333: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            334: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            335: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            336: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            337: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            338: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            339: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            340: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            341: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            342: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            343: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            344: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            345: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            346: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            347: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            348: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            349: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            350: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            351: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            352: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            353: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            354: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            355: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            356: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            357: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            358: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            359: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            360: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            361: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            362: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            363: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            364: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            365: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            366: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            367: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            368: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            369: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            370: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            371: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            372: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            373: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            374: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            375: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            376: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            377: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            378: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            379: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            380: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            381: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            382: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            383: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            384: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            385: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            386: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            387: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            388: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            389: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            390: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            391: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            392: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            393: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            394: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            395: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            396: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            397: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            398: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            399: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            400: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            401: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            402: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            403: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            404: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            405: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            406: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            407: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            408: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            409: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            410: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            411: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            412: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            413: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            414: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            415: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            416: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            417: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            418: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            419: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            420: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            421: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            422: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            423: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            424: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            425: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            426: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            427: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            428: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            429: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            430: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            431: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            432: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            433: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            434: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            435: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            436: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            437: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            438: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            439: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            440: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            441: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            442: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            443: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            444: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            445: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            446: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            447: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            448: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            449: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            450: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            451: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            452: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            453: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            454: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            455: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            456: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            457: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            458: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            459: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            460: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            461: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            462: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            463: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            464: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            465: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            466: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            467: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            468: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            469: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            470: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            471: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            472: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            473: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            474: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            475: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            476: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            477: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            478: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            479: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            480: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            481: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            482: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            483: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            484: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            485: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            486: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            487: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            488: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            489: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            490: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            491: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            492: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            493: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            494: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            495: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            496: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            497: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            498: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            499: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            500: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            501: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            502: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            503: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            504: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            505: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            506: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            507: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            508: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            509: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            510: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            511: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            512: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            513: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            514: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            515: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            516: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            517: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            518: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            519: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            520: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            521: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            522: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            523: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            524: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            525: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            526: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            527: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            528: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            529: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            530: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            531: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            532: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            533: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            534: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            535: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            536: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            537: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            538: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            539: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            540: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            541: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            542: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            543: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            544: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            545: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            546: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            547: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            548: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            549: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            550: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            551: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            552: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            553: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            554: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            555: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            556: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            557: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            558: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            559: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            560: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            561: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            562: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            563: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            564: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            565: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            566: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            567: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            568: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            569: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            570: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            571: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            572: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            573: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            574: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            575: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            576: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            577: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            578: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            579: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            580: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            581: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            582: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            583: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            584: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            585: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            586: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            587: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            588: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            589: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            590: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            591: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            592: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            593: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            594: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            595: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            596: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            597: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            598: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            599: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            600: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            601: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            602: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            603: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            604: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            605: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            606: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            607: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            608: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            609: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            610: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            611: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            612: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            613: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            614: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            615: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            616: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            617: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            618: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            619: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            620: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            621: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            622: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            623: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            624: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            625: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            626: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            627: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            628: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            629: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            630: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            631: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            632: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            633: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            634: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            635: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            636: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            637: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            638: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            639: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            640: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            641: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            642: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            643: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            644: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            645: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            646: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            647: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            648: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            649: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            650: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            651: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            652: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            653: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            654: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            655: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            656: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            657: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            658: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            659: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            660: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            661: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            662: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            663: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            664: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            665: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            666: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            667: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            668: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            669: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            670: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            671: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            672: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            673: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            674: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            675: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            676: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            677: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            678: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            679: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            680: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            681: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            682: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            683: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            684: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            685: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            686: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            687: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            688: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            689: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            690: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            691: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            692: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            693: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            694: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            695: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            696: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            697: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            698: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            699: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            700: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            701: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            702: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            703: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            704: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            705: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            706: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            707: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            708: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            709: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            710: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            711: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            712: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            713: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            714: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            715: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            716: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            717: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            718: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            719: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            720: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            721: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            722: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            723: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            724: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            725: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            726: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            727: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            728: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            729: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            730: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            731: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            732: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            733: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            734: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            735: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            736: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            737: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            738: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            739: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            740: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            741: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            742: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            743: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            744: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            745: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            746: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            747: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            748: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            749: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            750: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            751: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            752: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            753: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            754: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            755: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            756: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            757: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            758: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            759: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            760: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            761: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            762: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            763: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            764: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            765: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            766: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            767: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            768: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            769: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            770: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            771: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            772: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            773: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            774: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            775: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            776: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            777: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            778: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            779: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            780: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            781: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            782: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            783: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            784: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            785: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            786: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            787: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            788: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            789: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            790: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            791: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            792: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            793: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            794: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_0A5B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            2: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            3: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            4: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            5: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            6: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            7: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            8: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            9: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            10: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            11: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            12: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            13: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            14: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            15: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            16: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            17: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            18: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            19: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            20: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            21: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            22: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            23: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            24: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            25: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            26: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            27: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            28: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            29: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            30: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            31: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            32: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            33: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            34: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            35: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            36: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            37: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            38: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            39: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            40: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            41: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            42: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            43: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_0A3B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            1: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            2: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            3: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            4: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            5: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            6: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            7: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            8: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            9: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            10: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            11: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            12: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            13: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            14: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            15: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            16: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            17: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            18: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            19: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            20: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            21: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            22: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            23: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            24: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            25: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            26: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            27: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            28: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            29: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            30: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            31: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            32: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            33: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            34: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            35: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            36: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            37: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            38: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            39: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            40: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            41: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            42: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            43: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            44: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            45: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            46: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            47: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            48: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            49: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            50: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            51: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            52: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            53: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            54: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            55: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            56: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            57: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            58: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            59: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            60: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            61: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            62: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            63: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            64: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            65: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            66: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            67: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            68: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            69: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            70: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            71: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            72: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            73: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            74: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            75: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            76: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            77: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            78: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            79: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            80: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            81: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            82: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            83: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            84: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            85: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            86: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            87: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            88: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            89: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            90: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            91: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            92: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            93: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            94: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            95: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            96: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            97: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            98: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            99: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            100: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            101: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            102: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            103: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            104: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            105: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            106: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            107: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            108: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            109: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            110: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            111: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            112: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            113: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            114: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            115: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            116: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            117: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            118: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            119: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            120: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            121: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            122: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            123: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            124: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            125: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            126: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            127: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            128: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            129: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            130: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            131: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            132: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            133: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            134: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            135: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            136: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            137: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            138: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            139: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            140: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            141: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            142: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            143: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            144: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            145: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            146: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            147: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            148: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            149: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            150: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            151: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            152: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            153: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            154: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            155: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            156: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            157: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            158: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            159: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            160: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            161: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            162: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            163: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            164: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            165: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            166: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            167: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            168: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            169: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            170: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            171: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            172: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            173: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            174: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            175: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            176: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            177: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            178: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            179: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            180: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            181: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            182: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            183: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            184: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            185: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            186: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            187: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            188: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            189: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            190: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            191: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            192: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            193: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            194: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            195: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            196: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            197: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            198: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            199: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            200: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            201: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            202: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            203: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            204: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            205: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            206: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            207: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            208: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            209: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            210: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            211: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            212: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            213: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            214: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            215: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            216: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            217: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            218: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            219: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            220: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            221: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            222: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            223: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            224: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            225: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            226: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            227: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            228: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            229: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            230: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            231: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            232: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            233: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            234: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            235: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            236: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            237: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            238: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            239: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            240: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            241: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            242: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            243: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            244: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            245: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            246: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            247: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            248: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            249: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            250: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            251: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            252: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            253: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            254: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            255: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            256: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            257: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            258: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            259: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            260: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            261: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            262: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            263: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            264: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            265: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            266: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            267: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            268: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            269: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            270: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            271: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            272: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            273: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            274: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            275: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            276: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            277: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            278: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            279: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            280: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            281: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            282: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            283: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            284: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            285: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            286: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            287: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            288: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            289: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            290: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            291: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            292: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            293: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            294: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            295: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            296: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            297: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            298: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            299: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            300: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            301: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            302: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            303: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            304: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            305: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            306: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            307: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            308: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            309: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            310: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            311: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            312: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            313: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            314: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            315: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            316: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            317: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            318: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            319: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            320: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            321: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            322: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            323: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            324: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            325: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            326: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            327: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            328: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            329: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            330: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            331: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            332: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            333: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            334: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            335: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            336: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            337: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            338: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            339: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            340: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            341: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            342: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            343: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            344: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            345: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            346: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            347: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            348: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            349: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            350: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            351: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            352: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            353: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            354: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            355: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            356: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            357: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            358: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            359: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            360: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            361: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            362: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            363: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            364: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            365: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            366: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            367: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            368: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            369: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            370: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            371: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            372: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            373: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            374: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            375: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            376: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            377: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            378: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            379: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            380: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            381: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            382: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            383: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            384: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            385: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            386: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            387: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            388: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            389: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            390: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            391: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            392: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            393: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            394: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            395: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            396: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            397: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            398: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            399: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            400: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            401: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            402: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            403: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            404: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            405: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            406: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            407: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            408: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            409: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            410: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            411: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            412: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            413: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            414: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            415: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            416: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            417: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            418: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            419: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            420: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            421: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            422: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            423: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            424: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            425: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            426: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            427: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            428: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            429: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            430: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            431: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            432: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            433: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            434: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            435: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            436: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            437: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            438: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            439: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            440: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            441: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            442: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            443: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            444: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            445: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            446: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            447: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            448: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            449: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            450: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            451: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            452: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            453: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            454: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            455: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            456: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            457: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            458: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            459: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            460: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            461: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            462: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            463: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            464: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            465: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            466: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            467: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            468: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            469: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            470: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            471: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            472: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            473: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            474: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            475: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            476: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            477: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            478: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            479: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            480: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            481: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            482: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            483: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            484: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            485: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            486: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            487: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            488: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            489: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            490: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            491: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            492: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            493: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            494: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            495: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            496: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            497: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            498: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            499: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            500: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            501: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            502: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            503: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            504: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            505: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            506: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            507: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            508: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            509: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            510: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            511: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            512: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            513: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            514: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            515: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            516: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            517: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            518: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            519: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            520: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            521: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            522: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            523: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            524: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            525: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            526: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            527: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            528: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            529: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            530: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            531: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            532: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            533: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            534: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            535: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            536: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            537: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            538: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            539: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            540: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            541: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            542: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            543: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            544: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            545: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            546: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            547: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            548: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            549: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            550: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            551: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            552: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            553: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            554: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            555: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            556: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            557: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            558: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            559: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            560: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            561: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            562: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            563: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            564: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            565: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            566: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            567: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            568: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            569: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            570: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            571: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            572: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            573: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            574: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            575: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            576: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            577: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            578: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            579: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            580: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            581: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            582: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            583: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            584: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            585: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            586: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            587: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            588: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            589: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            590: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            591: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            592: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            593: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            594: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            595: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            596: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            597: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            598: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            599: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            600: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            601: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            602: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            603: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            604: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            605: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            606: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            607: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            608: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            609: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            610: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            611: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            612: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            613: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            614: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            615: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            616: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            617: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            618: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            619: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            620: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            621: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            622: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            623: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            624: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            625: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            626: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            627: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            628: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            629: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            630: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            631: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            632: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            633: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            634: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            635: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            636: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            637: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            638: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            639: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            640: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            641: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            642: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            643: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            644: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            645: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            646: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            647: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            648: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            649: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            650: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            651: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            652: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            653: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            654: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            655: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            656: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            657: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            658: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            659: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            660: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            661: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            662: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            663: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            664: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            665: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            666: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            667: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            668: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            669: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            670: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            671: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            672: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            673: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            674: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            675: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            676: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            677: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            678: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            679: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            680: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            681: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            682: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            683: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            684: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            685: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            686: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            687: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            688: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            689: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            690: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            691: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            692: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            693: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            694: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            695: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            696: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            697: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            698: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            699: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            700: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            701: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            702: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            703: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            704: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            705: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            706: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            707: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            708: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            709: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            710: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            711: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            712: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            713: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            714: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            715: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            716: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            717: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            718: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            719: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            720: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            721: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            722: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            723: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            724: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            725: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            726: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            727: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            728: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            729: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            730: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            731: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            732: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            733: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            734: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            735: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            736: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            737: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            738: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            739: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            740: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            741: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            742: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            743: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            744: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            745: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            746: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            747: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            748: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            749: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            750: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            751: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            752: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            753: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            754: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            755: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            756: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            757: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            758: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            759: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            760: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            761: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            762: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            763: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            764: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            765: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            766: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            767: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            768: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            769: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            770: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            771: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            772: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            773: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            774: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            775: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            776: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            777: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            778: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            779: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            780: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            781: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            782: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            783: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            784: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            785: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            786: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            787: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            788: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            789: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            790: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            791: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            792: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            793: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            794: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            795: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            796: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            797: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            798: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            799: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            800: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            801: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            802: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            803: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            804: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            805: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            806: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            807: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            808: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            809: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            810: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            811: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            812: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            813: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            814: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            815: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            816: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            817: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            818: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            819: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            820: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            821: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            822: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            823: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            824: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            825: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            826: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            827: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            828: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            829: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            830: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            831: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            832: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            833: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            834: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            835: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            836: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            837: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            838: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            839: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            840: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            841: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            842: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            843: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            844: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            845: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            846: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            847: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            848: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            849: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            850: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            851: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            852: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            853: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            854: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            855: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            856: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            857: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            858: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            859: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            860: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            861: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            862: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            863: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            864: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            865: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            866: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            867: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            868: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            869: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            870: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            871: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            872: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            873: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            874: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            875: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            876: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            877: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            878: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            879: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            880: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            881: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            882: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            883: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            884: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            885: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            886: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            887: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            888: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            889: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            890: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            891: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            892: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            893: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            894: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            895: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            896: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            897: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            898: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            899: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            900: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            901: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            902: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            903: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            904: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            905: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            906: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            907: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            908: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            909: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            910: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            911: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            912: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            913: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            914: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            915: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            916: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            917: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            918: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            919: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            920: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            921: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            922: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            923: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            924: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            925: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            926: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            927: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            928: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            929: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            930: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            931: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            932: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            933: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            934: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            935: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            936: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            937: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            938: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            939: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            940: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            941: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            942: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            943: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            944: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            945: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            946: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            947: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            948: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            949: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            950: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            951: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            952: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            953: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            954: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            955: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            956: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            957: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            958: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            959: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            960: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            961: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            962: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            963: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            964: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            965: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            966: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            967: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            968: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            969: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            970: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            971: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            972: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            973: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            974: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            975: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            976: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            977: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            978: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            979: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            980: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            981: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            982: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            983: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            984: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            985: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            986: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            987: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            988: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            989: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            990: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            991: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            992: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            993: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            994: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            995: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            996: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            997: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            998: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            999: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1000: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1001: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1002: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1003: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1004: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1005: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1006: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1007: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1008: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1009: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1010: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1011: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1012: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1013: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1014: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1015: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1016: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1017: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1018: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1019: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1020: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1021: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1022: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1023: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1024: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1025: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1026: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1027: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1028: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1029: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1030: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1031: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1032: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1033: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1034: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1035: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1036: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1037: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1038: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1039: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1040: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1041: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1042: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1043: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1044: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1045: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1046: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1047: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1048: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1049: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1050: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1051: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1052: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1053: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1054: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1055: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1056: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1057: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1058: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1059: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1060: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1061: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1062: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1063: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1064: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1065: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1066: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1067: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1068: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1069: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1070: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1071: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1072: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1073: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1074: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1075: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1076: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1077: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1078: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1079: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1080: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1081: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1082: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1083: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1084: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1085: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1086: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1087: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1088: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1089: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1090: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1091: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1092: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1093: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1094: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1095: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1096: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1097: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1098: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1099: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1100: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1101: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1102: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1103: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1104: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1105: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1106: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1107: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1108: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1109: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1110: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1111: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1112: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1113: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1114: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1115: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1116: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1117: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1118: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1119: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1120: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1121: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1122: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1123: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1124: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1125: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1126: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1127: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1128: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1129: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1130: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1131: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1132: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1133: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1134: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1135: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1136: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1137: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1138: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1139: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1140: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1141: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1142: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1143: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1144: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1145: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1146: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1147: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1148: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1149: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1150: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1151: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1152: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1153: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1154: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1155: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1156: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1157: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1158: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1159: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1160: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1161: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1162: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1163: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1164: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1165: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1166: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1167: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1168: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1169: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1170: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1171: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1172: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1173: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1174: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1175: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1176: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1177: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1178: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1179: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1180: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1181: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1182: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1183: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1184: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1185: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1186: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1187: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1188: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1189: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1190: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1191: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1192: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1193: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1194: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1195: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1196: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1197: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1198: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1199: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1200: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1201: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1202: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1203: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1204: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1205: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1206: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1207: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1208: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1209: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1210: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1211: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1212: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1213: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1214: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1215: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1216: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1217: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1218: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1219: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1220: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1221: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1222: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1223: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1224: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1225: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1226: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1227: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1228: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1229: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1230: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1231: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1232: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1233: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1234: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1235: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1236: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1237: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1238: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1239: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1240: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1241: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1242: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1243: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1244: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1245: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1246: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1247: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1248: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1249: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1250: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1251: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1252: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1253: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1254: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1255: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1256: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1257: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1258: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1259: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1260: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1261: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1262: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1263: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1264: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1265: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1266: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1267: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1268: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1269: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1270: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1271: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1272: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1273: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1274: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1275: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1276: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1277: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1278: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1279: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1280: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1281: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1282: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1283: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1284: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1285: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1286: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1287: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1288: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1289: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1290: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1291: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1292: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1293: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1294: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1295: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1296: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1297: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1298: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1299: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1300: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1301: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1302: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1303: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1304: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1305: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1306: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1307: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1308: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1309: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1310: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1311: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1312: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1313: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1314: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1315: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1316: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1317: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1318: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1319: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1320: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1321: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1322: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1323: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1324: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1325: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1326: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1327: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1328: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1329: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1330: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1331: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1332: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1333: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1334: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1335: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1336: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1337: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1338: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1339: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1340: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1341: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1342: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1343: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1344: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1345: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1346: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1347: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1348: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1349: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1350: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1351: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1352: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1353: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1354: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1355: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1356: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1357: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1358: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1359: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1360: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1361: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1362: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1363: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1364: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1365: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1366: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1367: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1368: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1369: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1370: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1371: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1372: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1373: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1374: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1375: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1376: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1377: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1378: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1379: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1380: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1381: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1382: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1383: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1384: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1385: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1386: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1387: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1388: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1389: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1390: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1391: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1392: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1393: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1394: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1395: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1396: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1397: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1398: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1399: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1400: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1401: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1402: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1403: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1404: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1405: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1406: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1407: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1408: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1409: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1410: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1411: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1412: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1413: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1414: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1415: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1416: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1417: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1418: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1419: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1420: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1421: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1422: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1423: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1424: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1425: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1426: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1427: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1428: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1429: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1430: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1431: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1432: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1433: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1434: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1435: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1436: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1437: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1438: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1439: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1440: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1441: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1442: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1443: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1444: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1445: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1446: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1447: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1448: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1449: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1450: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1451: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1452: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1453: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1454: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1455: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1456: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1457: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1458: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1459: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1460: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1461: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1462: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1463: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1464: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1465: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1466: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1467: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1468: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1469: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1470: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1471: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1472: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1473: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1474: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1475: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1476: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1477: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1478: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1479: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1480: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1481: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1482: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1483: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1484: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1485: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1486: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1487: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1488: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1489: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1490: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1491: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1492: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1493: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1494: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1495: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1496: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1497: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1498: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1499: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1500: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1501: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1502: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1503: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1504: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1505: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1506: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1507: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1508: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1509: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1510: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1511: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1512: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1513: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1514: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1515: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            1516: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1517: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1518: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1519: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1520: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1521: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1522: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1523: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1524: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1525: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1526: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1527: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1528: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1529: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1530: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1531: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1532: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1533: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1534: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1535: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1536: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1537: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1538: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1539: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1540: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1541: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1542: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1543: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1544: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1545: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1546: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1547: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1548: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1549: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1550: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1551: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1552: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1553: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1554: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1555: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1556: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1557: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1558: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1559: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1560: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1561: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1562: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1563: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1564: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1565: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1566: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1567: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1568: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1569: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            1570: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1571: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            1572: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1573: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            1574: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1575: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            1576: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1577: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1578: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1579: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            1580: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            1581: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            1582: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1583: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1584: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1585: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1586: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1587: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1588: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1589: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1590: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1591: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1592: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1593: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1594: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1595: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1596: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1597: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1598: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1599: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1600: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1601: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1602: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1603: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1604: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1605: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1606: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1607: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1608: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1609: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1610: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1611: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1612: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1613: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1614: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1615: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1616: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1617: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1618: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1619: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1620: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1621: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1622: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1623: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1624: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1625: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1626: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1627: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1628: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1629: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1630: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1631: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1632: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1633: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1634: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1635: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1636: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1637: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1638: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1639: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1640: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1641: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1642: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1643: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1644: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1645: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1646: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1647: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1648: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1649: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1650: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1651: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1652: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1653: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1654: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1655: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1656: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1657: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1658: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1659: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1660: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1661: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1662: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1663: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1664: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1665: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1666: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1667: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1668: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1669: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1670: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1671: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1672: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1673: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1674: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1675: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1676: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1677: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1678: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1679: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1680: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1681: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1682: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1683: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1684: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1685: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1686: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1687: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1688: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1689: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1690: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1691: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1692: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1693: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1694: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1695: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1696: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1697: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1698: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1699: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1700: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1701: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1702: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1703: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1704: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1705: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1706: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1707: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1708: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1709: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1710: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1711: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1712: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1713: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1714: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1715: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1716: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1717: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1718: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1719: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1720: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1721: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1722: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1723: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1724: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1725: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1726: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1727: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1728: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1729: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1730: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1731: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1732: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1733: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1734: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1735: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1736: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1737: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1738: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1739: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1740: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1741: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1742: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1743: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1744: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1745: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1746: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1747: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1748: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1749: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1750: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1751: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1752: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1753: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1754: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1755: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1756: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1757: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1758: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1759: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1760: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1761: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1762: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1763: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1764: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1765: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1766: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1767: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1768: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1769: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1770: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            1771: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            1772: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1773: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1774: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1775: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1776: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1777: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1778: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1779: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1780: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1781: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1782: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1783: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1784: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1785: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1786: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1787: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1788: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1789: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1790: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1791: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1792: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1793: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1794: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1795: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1796: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1797: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1798: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1799: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1800: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1801: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1802: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1803: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1804: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1805: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1806: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1807: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1808: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1809: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1810: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1811: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1812: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1813: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1814: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1815: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1816: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1817: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1818: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1819: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1820: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1821: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1822: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            1823: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1824: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1825: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            1826: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            1827: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            1828: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            1829: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            1830: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            1831: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            1832: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            1833: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            1834: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            1835: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            1836: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            1837: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            1838: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1839: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1840: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1841: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1842: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1843: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1844: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1845: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1846: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1847: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1848: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1849: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1850: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1851: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1852: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1853: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1854: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1855: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1856: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1857: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1858: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1859: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1860: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1861: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1862: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1863: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1864: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1865: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1866: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1867: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1868: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1869: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1870: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1871: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1872: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1873: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1874: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1875: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1876: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1877: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1878: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1879: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1880: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1881: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1882: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1883: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1884: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1885: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1886: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1887: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1888: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1889: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1890: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1891: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1892: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1893: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1894: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1895: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1896: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1897: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1898: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            1899: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1900: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1901: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            1902: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1903: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1904: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1905: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1906: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1907: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1908: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            1909: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            1910: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            1911: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            1912: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            1913: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            1914: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            1915: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            1916: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            1917: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            1918: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            1919: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        STATE_0A2B: case (cnt)
            0: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            1: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            2: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            3: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            4: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            5: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            6: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            7: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            8: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            9: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            10: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            11: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            12: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            13: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            14: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            15: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            16: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            17: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            18: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            19: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            20: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            21: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            22: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            23: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            24: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            25: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            26: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            27: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            28: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            29: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            30: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            31: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            32: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            33: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            34: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            35: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            36: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            37: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            38: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            39: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            40: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            41: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            42: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            43: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            44: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            45: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            46: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            47: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            48: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            49: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            50: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            51: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            52: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            53: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            54: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            55: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            56: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            57: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            58: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            59: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            60: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            61: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            62: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            63: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            64: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            65: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            66: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            67: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            68: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            69: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            70: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            71: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            72: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            73: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            74: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            75: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            76: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            77: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            78: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            79: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            80: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            81: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            82: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            83: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            84: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            85: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            86: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            87: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            88: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            89: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            90: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            91: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            92: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            93: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            94: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            95: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            96: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            97: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            98: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            99: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            100: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            101: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            102: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            103: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            104: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            105: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            106: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            107: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            108: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            109: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            110: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            111: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            112: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            113: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            114: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            115: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            116: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            117: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            118: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            119: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            120: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            121: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            122: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            123: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            124: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            125: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            126: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            127: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            128: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            129: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            130: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            131: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            132: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            133: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            134: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            135: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            136: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            137: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            138: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            139: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            140: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            141: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            142: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            143: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            144: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            145: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            146: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            147: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            148: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            149: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            150: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            151: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            152: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            153: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            154: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            155: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            156: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            157: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            158: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            159: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            160: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            161: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            162: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            163: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            164: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            165: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            166: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            167: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            168: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            169: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            170: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            171: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            172: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            173: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            174: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            175: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            176: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            177: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            178: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            179: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            180: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            181: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            182: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            183: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            184: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            185: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            186: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            187: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            188: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            189: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            190: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            191: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            192: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            193: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            194: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            195: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            196: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            197: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            198: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            199: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            200: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            201: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            202: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            203: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            204: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            205: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            206: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            207: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            208: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            209: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            210: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            211: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            212: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            213: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            214: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            215: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            216: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            217: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            218: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            219: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            220: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            221: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            222: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            223: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            224: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            225: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            226: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            227: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            228: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            229: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            230: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            231: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            232: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            233: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            234: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            235: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            236: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            237: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            238: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            239: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            240: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            241: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            242: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            243: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            244: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            245: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            246: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            247: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            248: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            249: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            250: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            251: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            252: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            253: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            254: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            255: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            256: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            257: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            258: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            259: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            260: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            261: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            262: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            263: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            264: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            265: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            266: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            267: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            268: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            269: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            270: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            271: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            272: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            273: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            274: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            275: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            276: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            277: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            278: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            279: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            280: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            281: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            282: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            283: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            284: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            285: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            286: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            287: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            288: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            289: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            290: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            291: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            292: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            293: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            294: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            295: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            296: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            297: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            298: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            299: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            300: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            301: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            302: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            303: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            304: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            305: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            306: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            307: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            308: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            309: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            310: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            311: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            312: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            313: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            314: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            315: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            316: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            317: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            318: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            319: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            320: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            321: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            322: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            323: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            324: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            325: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            326: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            327: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            328: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            329: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            330: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            331: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            332: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            333: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            334: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            335: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            336: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            337: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            338: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            339: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            340: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            341: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            342: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            343: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            344: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            345: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            346: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            347: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            348: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            349: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            350: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            351: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            352: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            353: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            354: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            355: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            356: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            357: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            358: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            359: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            360: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            361: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            362: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            363: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            364: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            365: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            366: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            367: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            368: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            369: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            370: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            371: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            372: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            373: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            374: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            375: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            376: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            377: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            378: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            379: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            380: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            381: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            382: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            383: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            384: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            385: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            386: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            387: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            388: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            389: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            390: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            391: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            392: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            393: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            394: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            395: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            396: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            397: begin perm_arr[0]<=reorder_arr[5];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            398: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            399: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            400: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            401: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            402: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            403: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            404: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            405: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            406: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            407: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            408: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            409: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            410: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            411: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            412: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            413: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            414: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            415: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            416: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            417: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            418: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            419: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            420: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            421: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            422: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            423: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            424: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            425: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            426: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            427: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            428: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            429: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            430: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            431: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            432: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            433: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            434: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            435: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            436: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            437: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            438: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            439: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            440: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            441: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            442: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            443: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            444: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            445: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            446: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            447: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            448: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            449: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            450: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            451: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            452: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            453: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            454: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            455: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            456: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            457: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            458: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            459: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            460: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            461: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            462: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            463: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            464: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            465: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            466: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            467: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            468: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            469: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            470: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            471: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            472: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            473: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            474: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            475: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            476: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            477: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            478: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            479: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            480: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            481: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            482: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            483: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            484: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            485: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            486: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            487: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            488: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            489: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            490: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            491: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            492: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            493: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            494: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            495: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            496: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            497: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            498: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            499: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            500: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            501: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            502: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            503: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            504: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            505: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            506: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            507: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            508: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            509: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            510: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            511: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            512: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            513: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            514: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            515: begin perm_arr[0]<=reorder_arr[3];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            516: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            517: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            518: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            519: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            520: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            521: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            522: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            523: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            524: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            525: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            526: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            527: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            528: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            529: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            530: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            531: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            532: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            533: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            534: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            535: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            536: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            537: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            538: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            539: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            540: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            541: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            542: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            543: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            544: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            545: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            546: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            547: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            548: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            549: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            550: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            551: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            552: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            553: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            554: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            555: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            556: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            557: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            558: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            559: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            560: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            561: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            562: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            563: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            564: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            565: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            566: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            567: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            568: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            569: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            570: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            571: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            572: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            573: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            574: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            575: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            576: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            577: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            578: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            579: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            580: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            581: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            582: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            583: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            584: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            585: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            586: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            587: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            588: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            589: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            590: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            591: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            592: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            593: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            594: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[4];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            595: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            596: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            597: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            598: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            599: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            600: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            601: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            602: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            603: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            604: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            605: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            606: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            607: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            608: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            609: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            610: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            611: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            612: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            613: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            614: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            615: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            616: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            617: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            618: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            619: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[7]; end
            620: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            621: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            622: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            623: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            624: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            625: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            626: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            627: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            628: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            629: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            630: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            631: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            632: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            633: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            634: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            635: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            636: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            637: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            638: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            639: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            640: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            641: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            642: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            643: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            644: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            645: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            646: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            647: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            648: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            649: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            650: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            651: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            652: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            653: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            654: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            655: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            656: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            657: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            658: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            659: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            660: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            661: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            662: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            663: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            664: begin perm_arr[0]<=reorder_arr[1];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            665: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            666: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            667: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            668: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            669: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            670: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            671: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            672: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            673: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            674: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            675: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            676: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            677: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            678: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            679: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            680: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            681: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            682: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            683: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            684: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            685: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            686: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            687: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            688: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            689: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            690: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            691: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            692: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            693: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[1]; end
            694: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[2]; end
            695: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[3]; end
            696: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            697: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[0]; end
            698: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[2]; end
            699: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[3]; end
            700: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            701: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[0]; end
            702: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[1]; end
            703: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[3]; end
            704: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            705: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            706: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[0]; end
            707: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[1]; end
            708: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[2]; end
            709: begin perm_arr[0]<=reorder_arr[6];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[3]; end
            710: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            711: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            712: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            713: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            714: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            715: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            716: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            717: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            718: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            719: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            720: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            721: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            722: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            723: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[4];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            724: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            725: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            726: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            727: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            728: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            729: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            730: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[6]; end
            731: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            732: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            733: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            734: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            735: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            736: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            737: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            738: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            739: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            740: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            741: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[6]; end
            742: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[6]; end
            743: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[4];perm_arr[4]<=reorder_arr[5]; end
            744: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            745: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            746: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[6]; end
            747: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[0];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            748: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[0]; end
            749: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[1]; end
            750: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[2]; end
            751: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[5];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[3]; end
            752: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            753: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            754: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            755: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[1];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            756: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            757: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[3];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            758: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[7]; end
            759: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[7]; end
            760: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[6]; end
            761: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[7]; end
            762: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[7]; end
            763: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[0]; end
            764: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[1]; end
            765: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[2]; end
            766: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[5];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[3]; end
            767: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[7]; end
            768: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[0];perm_arr[4]<=reorder_arr[5]; end
            769: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[6];perm_arr[3]<=reorder_arr[7];perm_arr[4]<=reorder_arr[5]; end
            770: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[1];perm_arr[4]<=reorder_arr[5]; end
            771: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[2];perm_arr[4]<=reorder_arr[5]; end
            772: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[0]; end
            773: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[1]; end
            774: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[2]; end
            775: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[6];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[3]; end
            776: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            777: begin perm_arr[0]<=reorder_arr[2];perm_arr[1]<=reorder_arr[3];perm_arr[2]<=reorder_arr[7];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            778: begin perm_arr[0]<=reorder_arr[7];perm_arr[1]<=reorder_arr[2];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[6];perm_arr[4]<=reorder_arr[5]; end
            779: begin perm_arr[0]<=reorder_arr[4];perm_arr[1]<=reorder_arr[7];perm_arr[2]<=reorder_arr[0];perm_arr[3]<=reorder_arr[5];perm_arr[4]<=reorder_arr[6]; end
            default: begin perm_arr[0]<=0;perm_arr[1]<=0;perm_arr[2]<=0;perm_arr[3]<=0;perm_arr[4]<=0; end
        endcase
        default: begin
            perm_arr[0] <= 0;
            perm_arr[1] <= 0;
            perm_arr[2] <= 0;
            perm_arr[3] <= 0;
            perm_arr[4] <= 0;
        end
    endcase
end

always @(posedge clk or negedge rst_n) begin // calculate the weighted sum
    if (!rst_n) begin
        weighted_sum <= 0;
        weighted_sum_2 <= 0;
        bwnc <= 0;
        prev_perm_arr[0] <= 0;
        prev_perm_arr[1] <= 0;
        prev_perm_arr[2] <= 0;
        prev_perm_arr[3] <= 0;
        prev_perm_arr[4] <= 0;
    end
    else
    case (current_state)
        STATE_5A0B, STATE_4A0B, STATE_3A2B, STATE_3A1B, STATE_3A0B,
        STATE_2A2B, STATE_2A3B, STATE_2A1B, STATE_2A0B, STATE_1A4B,
        STATE_1A3B, STATE_1A2B, STATE_1A1B, STATE_0A4B, STATE_0A5B,
        STATE_0A3B, STATE_0A2B: begin 
            weighted_sum <= (weight_arr[0]*perm_arr[0]) + (weight_arr[1]*perm_arr[1]) + (weight_arr[2]*perm_arr[2]) + (weight_arr[3]*perm_arr[3]) + (weight_arr[4]*perm_arr[4]);
            weighted_sum_2 <= (16*perm_arr[0]) + (8*perm_arr[1]) + (4*perm_arr[2]) + (2*perm_arr[3]) + (1*perm_arr[4]);
            bwnc <= ~{perm_arr[0],perm_arr[1],perm_arr[2],perm_arr[3],perm_arr[4]};
            prev_perm_arr[0] <= perm_arr[0];
            prev_perm_arr[1] <= perm_arr[1];
            prev_perm_arr[2] <= perm_arr[2];
            prev_perm_arr[3] <= perm_arr[3];
            prev_perm_arr[4] <= perm_arr[4];    
        end
        default: begin
            weighted_sum <= 0;
            weighted_sum_2 <= 0;
            bwnc <= 0;
            prev_perm_arr[0] <= 0;
            prev_perm_arr[1] <= 0;
            prev_perm_arr[2] <= 0;
            prev_perm_arr[3] <= 0;
            prev_perm_arr[4] <= 0;
        end
    endcase
end

always @(posedge clk or negedge rst_n) begin // update the reuslt based on weighted sum
    if (!rst_n) begin
        max_weighted_sum <= 0;
        max_weighted_sum_2 <= 0;
        max_bwnc <= 0;
        result_arr[0] <= 0;
        result_arr[1] <= 0;
        result_arr[2] <= 0;
        result_arr[3] <= 0;
        result_arr[4] <= 0;
    end
    else
    case (current_state)
        STATE_5A0B, STATE_4A0B, STATE_3A2B, STATE_3A1B, STATE_3A0B,
        STATE_2A2B, STATE_2A3B, STATE_2A1B, STATE_2A0B, STATE_1A4B,
        STATE_1A3B, STATE_1A2B, STATE_1A1B, STATE_0A4B, STATE_0A5B,
        STATE_0A3B, STATE_0A2B: begin
            if (weighted_sum > max_weighted_sum) begin
                // valid, update result
                max_weighted_sum <= weighted_sum;
                max_weighted_sum_2 <= weighted_sum_2;
                max_bwnc <= bwnc;
                result_arr[0] <= prev_perm_arr[0];
                result_arr[1] <= prev_perm_arr[1];
                result_arr[2] <= prev_perm_arr[2];
                result_arr[3] <= prev_perm_arr[3];
                result_arr[4] <= prev_perm_arr[4];
            end
            else if (weighted_sum == max_weighted_sum) begin
                if (weighted_sum_2 > max_weighted_sum_2) begin
                    // valid, update result
                    max_weighted_sum <= weighted_sum;
                    max_weighted_sum_2 <= weighted_sum_2;
                    max_bwnc <= bwnc;
                    result_arr[0] <= prev_perm_arr[0];
                    result_arr[1] <= prev_perm_arr[1];
                    result_arr[2] <= prev_perm_arr[2];
                    result_arr[3] <= prev_perm_arr[3];
                    result_arr[4] <= prev_perm_arr[4];
                end
                else if (weighted_sum_2 == max_weighted_sum_2) begin
                    if (bwnc > max_bwnc) begin
                        // valid, update result
                        max_weighted_sum <= weighted_sum;
                        max_weighted_sum_2 <= weighted_sum_2;
                        max_bwnc <= bwnc;
                        result_arr[0] <= prev_perm_arr[0];
                        result_arr[1] <= prev_perm_arr[1];
                        result_arr[2] <= prev_perm_arr[2];
                        result_arr[3] <= prev_perm_arr[3];
                        result_arr[4] <= prev_perm_arr[4];
                    end
                    else begin
                        // invalid, remain unchanged
                        max_weighted_sum <= max_weighted_sum;
                        max_weighted_sum_2 <= max_weighted_sum_2;
                        max_bwnc <= max_bwnc;
                        result_arr[0] <= result_arr[0];
                        result_arr[1] <= result_arr[1];
                        result_arr[2] <= result_arr[2];
                        result_arr[3] <= result_arr[3];
                        result_arr[4] <= result_arr[4];
                    end
                end
                else begin
                    // invalid, remain unchanged
                    max_weighted_sum <= max_weighted_sum;
                    max_weighted_sum_2 <= max_weighted_sum_2;
                    max_bwnc <= max_bwnc;
                    result_arr[0] <= result_arr[0];
                    result_arr[1] <= result_arr[1];
                    result_arr[2] <= result_arr[2];
                    result_arr[3] <= result_arr[3];
                    result_arr[4] <= result_arr[4];
                end
            end
            else begin
                // invalid, remain unchanged
                max_weighted_sum <= max_weighted_sum;
                max_weighted_sum_2 <= max_weighted_sum_2;
                max_bwnc <= max_bwnc;
                result_arr[0] <= result_arr[0];
                result_arr[1] <= result_arr[1];
                result_arr[2] <= result_arr[2];
                result_arr[3] <= result_arr[3];
                result_arr[4] <= result_arr[4];
            end
        end
        STATE_OUTPUT: begin // reamin unchanged
            max_weighted_sum <= max_weighted_sum;
            max_weighted_sum_2 <= max_weighted_sum_2;
            max_bwnc <= max_bwnc;
            result_arr[0] <= result_arr[0];
            result_arr[1] <= result_arr[1];
            result_arr[2] <= result_arr[2];
            result_arr[3] <= result_arr[3];
            result_arr[4] <= result_arr[4];
        end 
        default: begin // zeroed
            max_weighted_sum <= 0;
            max_weighted_sum_2 <= 0;
            max_bwnc <= 0;
            result_arr[0] <= 0;
            result_arr[1] <= 0;
            result_arr[2] <= 0;
            result_arr[3] <= 0;
            result_arr[4] <= 0;
        end
    endcase
end

// Output logic
always @(posedge clk or negedge rst_n) begin // output out_valid
    if (!rst_n)
        out_valid <= 0;
    else
    case (current_state)
        STATE_OUTPUT: out_valid <= 1;
        default: out_valid <= 0;
    endcase
end
always @(posedge clk or negedge rst_n) begin // output result
    if (!rst_n) result <= 0;
    else
    case (current_state)
        STATE_OUTPUT:
        case (cnt)
            0: result <= result_arr[0]; 
            1: result <= result_arr[1]; 
            2: result <= result_arr[2]; 
            3: result <= result_arr[3];
            default: result <= result_arr[4];
        endcase
        default: result <= 0; 
    endcase
end
always @(posedge clk or negedge rst_n) begin // output out_value
    if (!rst_n) out_value <= 0;
    else
    case (current_state)
        STATE_OUTPUT: out_value <= max_weighted_sum; 
        default: out_value <= 0;
    endcase
end

endmodule